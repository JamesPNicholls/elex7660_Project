module joy_code(
    
);
    
endmodule