module parsse_adc(
    port_list
);
    
endmodule