/*********************************************************************
*BankVault Module (Top-level heirarchy)
*
*Date: 2/25/2022
*
*Author: Mo Amirian, Clint Gaudet, James Nicholls
*
*Class: ELEX 7660 - Digital System Design
*
*Module Description: 
*	Top level Entity used to handle state machine and individual modules
*
*
*
**********************************************************************/

module bankVault ( output logic [3:0] kpc,  // column select, active-low
              (* altera_attribute = "-name WEAK_PULL_UP_RESISTOR ON" *)
              input logic  [3:0] kpr,  // rows, active-low w/ pull-ups
              output logic [7:0] leds, // active-low LED segments 
              output logic [3:0] ct,   // " digit enables
              input logic  reset_n, FPGA_CLK1_50 ) ;

	logic clk ;                  // 2kHz clock for keypad scanning
	logic kphit ;                // a key is pressed
	logic [3:0] num ;            // value of pressed key
	logic [3:0] digit = 4'b0;
	logic [7:0] count = 'b0;	//counter for determining which 8-segment led
	pll pll0 ( .inclk0(FPGA_CLK1_50), .c0(clk) ) ;
	
  // Probably need anothe module to handle what and when things are sent to the LEDs
	always_ff@(posedge clk) begin
		if (kphit == 1'b1) begin
			while (kphit == 1'b1)
			digit[count] <= 1'b1;
			if (count >= 3)
				count <= 0;
			else
				count <= count + 1'b1;
		end

	end
	//assign ct = { {2{1'b0}}, kphit, kphit} ;
	assign ct = {digit[3], digit[2], digit[1], digit[0]} ;
	

	// instantiate your modules here...
	decode7 decode7_0 (.num,.leds) ;
	kpdecode kpdecode_0 (.kpr, .kpc, .kphit, .num);
	colseq colseq_0 (.clk, .reset_n, .kpr, .kpc);

  logic [7:0] current_state;
  logic [7:0] next_state;
  
  // System States
  localparam 
    start_up  = 0x0,
    game_1    = 0x1,
    game_2    = 0x2
    game_3    = 0x3,
    victory   = 0x4;
    fubar     = 0x5; //error state if anything bad happens

  // Almost everything should be inside this case statement
  // This block will decide what is sent to the the LEDS/7segs/etc
  // Also handles where the ADC, and keypad inputs will go
  always_comb begin : state_logic
    current_state = next_state;
    case (current_state)
      
      default: begin
        ;
      end
    endcase

  end : state_logic

  end

  // Handles state change in reponse to state logic 
  always_ff @( posedge clk, negedge reset_n ) begin : state_handler

    if(current_state == start_up      && /* Other */) begin
      next_state == game_1;
    end

    else if(current_state == game_1    && /* Other */) begin
      next_state = game_2
    end      

    else if(current_state == game_2    && /* Other */) begin
      next_state = game_3
    end

    else if(current_state == game_3    && /* Other */) begin
      next_state = victory
    end

    else if(current_state == victory   && /* Other */) begin
      next_state = fubar
    end

    else begin // WHEN EVERYTHING GOES WRONG
      next_state = current_state;
    end

  end : state_handler
   
endmodule



// megafunction wizard: %ALTPLL%
// ...
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
// ...

module pll ( inclk0, c0);

        input     inclk0;
        output    c0;

        wire [0:0] sub_wire2 = 1'h0;
        wire [4:0] sub_wire3;
        wire  sub_wire0 = inclk0;
        wire [1:0] sub_wire1 = {sub_wire2, sub_wire0};
        wire [0:0] sub_wire4 = sub_wire3[0:0];
        wire  c0 = sub_wire4;

        altpll altpll_component ( .inclk (sub_wire1), .clk
          (sub_wire3), .activeclock (), .areset (1'b0), .clkbad
          (), .clkena ({6{1'b1}}), .clkloss (), .clkswitch
          (1'b0), .configupdate (1'b0), .enable0 (), .enable1 (),
          .extclk (), .extclkena ({4{1'b1}}), .fbin (1'b1),
          .fbmimicbidir (), .fbout (), .fref (), .icdrclk (),
          .locked (), .pfdena (1'b1), .phasecounterselect
          ({4{1'b1}}), .phasedone (), .phasestep (1'b1),
          .phaseupdown (1'b1), .pllena (1'b1), .scanaclr (1'b0),
          .scanclk (1'b0), .scanclkena (1'b1), .scandata (1'b0),
          .scandataout (), .scandone (), .scanread (1'b0),
          .scanwrite (1'b0), .sclkout0 (), .sclkout1 (),
          .vcooverrange (), .vcounderrange ());

        defparam
                altpll_component.bandwidth_type = "AUTO",
                altpll_component.clk0_divide_by = 25000,
                altpll_component.clk0_duty_cycle = 50,
                altpll_component.clk0_multiply_by = 1,
                altpll_component.clk0_phase_shift = "0",
                altpll_component.compensate_clock = "CLK0",
                altpll_component.inclk0_input_frequency = 20000,
                altpll_component.intended_device_family = "Cyclone IV E",
                altpll_component.lpm_hint = "CBX_MODULE_PREFIX=lab1clk",
                altpll_component.lpm_type = "altpll",
                altpll_component.operation_mode = "NORMAL",
                altpll_component.pll_type = "AUTO",
                altpll_component.port_activeclock = "PORT_UNUSED",
                altpll_component.port_areset = "PORT_UNUSED",
                altpll_component.port_clkbad0 = "PORT_UNUSED",
                altpll_component.port_clkbad1 = "PORT_UNUSED",
                altpll_component.port_clkloss = "PORT_UNUSED",
                altpll_component.port_clkswitch = "PORT_UNUSED",
                altpll_component.port_configupdate = "PORT_UNUSED",
                altpll_component.port_fbin = "PORT_UNUSED",
                altpll_component.port_inclk0 = "PORT_USED",
                altpll_component.port_inclk1 = "PORT_UNUSED",
                altpll_component.port_locked = "PORT_UNUSED",
                altpll_component.port_pfdena = "PORT_UNUSED",
                altpll_component.port_phasecounterselect = "PORT_UNUSED",
                altpll_component.port_phasedone = "PORT_UNUSED",
                altpll_component.port_phasestep = "PORT_UNUSED",
                altpll_component.port_phaseupdown = "PORT_UNUSED",
                altpll_component.port_pllena = "PORT_UNUSED",
                altpll_component.port_scanaclr = "PORT_UNUSED",
                altpll_component.port_scanclk = "PORT_UNUSED",
                altpll_component.port_scanclkena = "PORT_UNUSED",
                altpll_component.port_scandata = "PORT_UNUSED",
                altpll_component.port_scandataout = "PORT_UNUSED",
                altpll_component.port_scandone = "PORT_UNUSED",
                altpll_component.port_scanread = "PORT_UNUSED",
                altpll_component.port_scanwrite = "PORT_UNUSED",
                altpll_component.port_clk0 = "PORT_USED",
                altpll_component.port_clk1 = "PORT_UNUSED",
                altpll_component.port_clk2 = "PORT_UNUSED",
                altpll_component.port_clk3 = "PORT_UNUSED",
                altpll_component.port_clk4 = "PORT_UNUSED",
                altpll_component.port_clk5 = "PORT_UNUSED",
                altpll_component.port_clkena0 = "PORT_UNUSED",
                altpll_component.port_clkena1 = "PORT_UNUSED",
                altpll_component.port_clkena2 = "PORT_UNUSED",
                altpll_component.port_clkena3 = "PORT_UNUSED",
                altpll_component.port_clkena4 = "PORT_UNUSED",
                altpll_component.port_clkena5 = "PORT_UNUSED",
                altpll_component.port_extclk0 = "PORT_UNUSED",
                altpll_component.port_extclk1 = "PORT_UNUSED",
                altpll_component.port_extclk2 = "PORT_UNUSED",
                altpll_component.port_extclk3 = "PORT_UNUSED",
                altpll_component.width_clock = 5;


endmodule

